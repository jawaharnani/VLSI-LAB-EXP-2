input d0,d1,d2,d3,d4,d5,d6,d7;

module encoder_8_to_3(a0,a1,a2,d0,d1,d2,d3,d4,d5,d6,d7); or g2(a1,d2,d3,d6,d7); or g3(a2,d4,d5,d6,d7);

output a0,a1,a2; or g1(a0,d1,d3,d5,d7);

endmodule
